module md5(
    input  clk,
    input  [0:63]  in_txt,
    output [0:127] hash,
    output [0:63]  out_txt  
);

localparam h0 = 32'h67452301;
localparam h1 = 32'hefcdab89;
localparam h2 = 32'h98badcfe;
localparam h3 = 32'h10325476;

reg [0:63] w, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63;
reg [0:31]                A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15, A16, A17, A18, A19, A20, A21, A22, A23, A24, A25, A26, A27, A28, A29, A30, A31, A32, A33, A34, A35, A36, A37, A38, A39, A40, A41, A42, A43, A44, A45, A46, A47, A48, A49, A50, A51, A52, A53, A54, A55, A56, A57, A58, A59, A60, A61, A62, A63;
reg [0:31]    B0, B1, B2, B3, B4, B5, B6, B7, B8, B9, B10, B11, B12, B13, B14, B15, B16, B17, B18, B19, B20, B21, B22, B23, B24, B25, B26, B27, B28, B29, B30, B31, B32, B33, B34, B35, B36, B37, B38, B39, B40, B41, B42, B43, B44, B45, B46, B47, B48, B49, B50, B51, B52, B53, B54, B55, B56, B57, B58, B59, B60, B61, B62, B63;
reg [0:31]        C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11, C12, C13, C14, C15, C16, C17, C18, C19, C20, C21, C22, C23, C24, C25, C26, C27, C28, C29, C30, C31, C32, C33, C34, C35, C36, C37, C38, C39, C40, C41, C42, C43, C44, C45, C46, C47, C48, C49, C50, C51, C52, C53, C54, C55, C56, C57, C58, C59, C60, C61, C62, C63;
reg [0:31]            D2, D3, D4, D5, D6, D7, D8, D9, D10, D11, D12, D13, D14, D15, D16, D17, D18, D19, D20, D21, D22, D23, D24, D25, D26, D27, D28, D29, D30, D31, D32, D33, D34, D35, D36, D37, D38, D39, D40, D41, D42, D43, D44, D45, D46, D47, D48, D49, D50, D51, D52, D53, D54, D55, D56, D57, D58, D59, D60, D61, D62, D63;

reg [0:127] hash_reg;
reg [0:63] out_reg;

assign hash = hash_reg;
assign out_txt = out_reg;

always @(posedge clk) begin
    w <= {in_txt[24+:8], in_txt[16+:8], in_txt[ 8+:8], in_txt[ 0+:8],
          in_txt[56+:8], in_txt[48+:8], in_txt[40+:8], in_txt[32+:8]};

    w0<=w;  w1<=w0; w2<=w1; w3<=w2; w4<=w3; w5<=w4; w6<=w5; w7<=w6; w8<=w7; w9 <=w8; w10<=w9;  w11<=w10; w12<=w11; w13<=w12; w14<=w13; w15<=w14; w16<=w15; w17<=w16; w18<=w17; w19<=w18; w20<=w19; w21<=w20; w22<=w21; w23<=w22; w24<=w23; w25<=w24; w26<=w25; w27<=w26; w28<=w27; w29<=w28; w30<=w29; w31<=w30; w32<=w31; w33<=w32; w34<=w33; w35<=w34; w36<=w35; w37<=w36; w38<=w37; w39<=w38; w40<=w39; w41<=w40; w42<=w41; w43<=w42; w44<=w43; w45<=w44; w46<=w45; w47<=w46; w48<=w47; w49<=w48; w50<=w49; w51<=w50; w52<=w51; w53<=w52; w54<=w53; w55<=w54; w56<=w55; w57<=w56; w58<=w57; w59<=w58; w60<=w59; w61<=w60; w62<=w61; w63<=w62;
                    A3<=D2; A4<=D3; A5<=D4; A6<=D5; A7<=D6; A8<=D7; A9<=D8; A10<=D9; A11<=D10; A12<=D11; A13<=D12; A14<=D13; A15<=D14; A16<=D15; A17<=D16; A18<=D17; A19<=D18; A20<=D19; A21<=D20; A22<=D21; A23<=D22; A24<=D23; A25<=D24; A26<=D25; A27<=D26; A28<=D27; A29<=D28; A30<=D29; A31<=D30; A32<=D31; A33<=D32; A34<=D33; A35<=D34; A36<=D35; A37<=D36; A38<=D37; A39<=D38; A40<=D39; A41<=D40; A42<=D41; A43<=D42; A44<=D43; A45<=D44; A46<=D45; A47<=D46; A48<=D47; A49<=D48; A50<=D49; A51<=D50; A52<=D51; A53<=D52; A54<=D53; A55<=D54; A56<=D55; A57<=D56; A58<=D57; A59<=D58; A60<=D59; A61<=D60; A62<=D61;
    C1<=B0; C2<=B1; C3<=B2; C4<=B3; C5<=B4; C6<=B5; C7<=B6; C8<=B7; C9<=B8; C10<=B9; C11<=B10; C12<=B11; C13<=B12; C14<=B13; C15<=B14; C16<=B15; C17<=B16; C18<=B17; C19<=B18; C20<=B19; C21<=B20; C22<=B21; C23<=B22; C24<=B23; C25<=B24; C26<=B25; C27<=B26; C28<=B27; C29<=B28; C30<=B29; C31<=B30; C32<=B31; C33<=B32; C34<=B33; C35<=B34; C36<=B35; C37<=B36; C38<=B37; C39<=B38; C40<=B39; C41<=B40; C42<=B41; C43<=B42; C44<=B43; C45<=B44; C46<=B45; C47<=B46; C48<=B47; C49<=B48; C50<=B49; C51<=B50; C52<=B51; C53<=B52; C54<=B53; C55<=B54; C56<=B55; C57<=B56; C58<=B57; C59<=B58; C60<=B59; C61<=B60; C62<=B61;
            D2<=C1; D3<=C2; D4<=C3; D5<=C4; D6<=C5; D7<=C6; D8<=C7; D9<=C8; D10<=C9; D11<=C10; D12<=C11; D13<=C12; D14<=C13; D15<=C14; D16<=C15; D17<=C16; D18<=C17; D19<=C18; D20<=C19; D21<=C20; D22<=C21; D23<=C22; D24<=C23; D25<=C24; D26<=C25; D27<=C26; D28<=C27; D29<=C28; D30<=C29; D31<=C30; D32<=C31; D33<=C32; D34<=C33; D35<=C34; D36<=C35; D37<=C36; D38<=C37; D39<=C38; D40<=C39; D41<=C40; D42<=C41; D43<=C42; D44<=C43; D45<=C44; D46<=C45; D47<=C46; D48<=C47; D49<=C48; D50<=C49; D51<=C50; D52<=C51; D53<=C52; D54<=C53; D55<=C54; D56<=C55; D57<=C56; D58<=C57; D59<=C58; D60<=C59; D61<=C60; D62<=C61;
    A63 <= D62 + h0;  C63 <= B62 + h2;  D63 <= C62 + h3;

    hash_reg <= {A63[24 +: 8], A63[16 +: 8], A63[ 8 +: 8], A63[ 0 +: 8],
                 B63[24 +: 8], B63[16 +: 8], B63[ 8 +: 8], B63[ 0 +: 8],
                 C63[24 +: 8], C63[16 +: 8], C63[ 8 +: 8], C63[ 0 +: 8],
                 D63[24 +: 8], D63[16 +: 8], D63[ 8 +: 8], D63[ 0 +: 8]};

    out_reg  <= {w63[24 +: 8], w63[16 +: 8], w63[ 8 +: 8], w63[ 0 +: 8],
                 w63[56 +: 8], w63[48 +: 8], w63[40 +: 8], w63[32 +: 8]};

    B0  <= (((32'hd76aa477                                     + w [0  +: 32]) <<  7)  |
            ((32'hd76aa478                                     + w [0  +: 32]) >> 25)) + h1;
    B1  <= (((32'hf8fa0bcc + ((B0 &h1 ) | ((~B0 )&h2 ))        + w0[32 +: 32]) << 12)  |
            ((32'hf8fa0bcc + ((B0 &h1 ) | ((~B0 )&h2 ))        + w0[32 +: 32]) >> 20)) + B0;
    B2  <= (((32'hbcdb4e59 + ((B1 &C1 ) | ((~B1 )&h1 ))                      ) << 17)  |
            ((32'hbcdb4e59 + ((B1 &C1 ) | ((~B1 )&h1 ))                      ) >> 15)) + B1;
    B3  <= (((32'hb18b7a77 + ((B2 &C2 ) | ((~B2 )&D2 ))                      ) << 22)  |
            ((32'hb18b7a77 + ((B2 &C2 ) | ((~B2 )&D2 ))                      ) >> 10)) + B2;
    B4  <= (((32'hf57c0faf + ((B3 &C3 ) | ((~B3 )&D3 )) + A3                 ) <<  7)  |
            ((32'hf57c0faf + ((B3 &C3 ) | ((~B3 )&D3 )) + A3                 ) >> 25)) + B3;
    B5  <= (((32'h4787c62a + ((B4 &C4 ) | ((~B4 )&D4 )) + A4                 ) << 12)  |
            ((32'h4787c62a + ((B4 &C4 ) | ((~B4 )&D4 )) + A4                 ) >> 20)) + B4;
    B6  <= (((32'ha8304613 + ((B5 &C5 ) | ((~B5 )&D5 )) + A5                 ) << 17)  |
            ((32'ha8304613 + ((B5 &C5 ) | ((~B5 )&D5 )) + A5                 ) >> 15)) + B5;
    B7  <= (((32'hfd469501 + ((B6 &C6 ) | ((~B6 )&D6 )) + A6                 ) << 22)  |
            ((32'hfd469501 + ((B6 &C6 ) | ((~B6 )&D6 )) + A6                 ) >> 10)) + B6;
    B8  <= (((32'h698098d8 + ((B7 &C7 ) | ((~B7 )&D7 )) + A7                 ) <<  7)  |
            ((32'h698098d8 + ((B7 &C7 ) | ((~B7 )&D7 )) + A7                 ) >> 25)) + B7;
    B9  <= (((32'h8b44f7af + ((B8 &C8 ) | ((~B8 )&D8 )) + A8                 ) << 12)  |
            ((32'h8b44f7af + ((B8 &C8 ) | ((~B8 )&D8 )) + A8                 ) >> 20)) + B8;
    B10 <= (((32'hffff5bb1 + ((B9 &C9 ) | ((~B9 )&D9 )) + A9                 ) << 17)  |
            ((32'hffff5bb1 + ((B9 &C9 ) | ((~B9 )&D9 )) + A9                 ) >> 15)) + B9;
    B11 <= (((32'h895cd7be + ((B10&C10) | ((~B10)&D10)) + A10                ) << 22)  |
            ((32'h895cd7be + ((B10&C10) | ((~B10)&D10)) + A10                ) >> 10)) + B10;
    B12 <= (((32'h6b901122 + ((B11&C11) | ((~B11)&D11)) + A11                ) <<  7)  |
            ((32'h6b901122 + ((B11&C11) | ((~B11)&D11)) + A11                ) >> 25)) + B11;
    B13 <= (((32'hfd987193 + ((B12&C12) | ((~B12)&D12)) + A12                ) << 12)  |
            ((32'hfd987193 + ((B12&C12) | ((~B12)&D12)) + A12                ) >> 20)) + B12;
    B14 <= (((32'ha67943ce + ((B13&C13) | ((~B13)&D13)) + A13                ) << 17)  |
            ((32'ha67943ce + ((B13&C13) | ((~B13)&D13)) + A13                ) >> 15)) + B13;
    B15 <= (((32'h49b40821 + ((B14&C14) | ((~B14)&D14)) + A14                ) << 22)  |
            ((32'h49b40821 + ((B14&C14) | ((~B14)&D14)) + A14                ) >> 10)) + B14;

    B16 <= (((32'hf61e2562 + ((D15&B15) | ((~D15)&C15)) + A15 + w15[32 +: 32]) <<  5)  |
            ((32'hf61e2562 + ((D15&B15) | ((~D15)&C15)) + A15 + w15[32 +: 32]) >> 27)) + B15;
    B17 <= (((32'hc040b340 + ((D16&B16) | ((~D16)&C16)) + A16                ) <<  9)  |
            ((32'hc040b340 + ((D16&B16) | ((~D16)&C16)) + A16                ) >> 23)) + B16;
    B18 <= (((32'h265e5a51 + ((D17&B17) | ((~D17)&C17)) + A17                ) << 14)  |
            ((32'h265e5a51 + ((D17&B17) | ((~D17)&C17)) + A17                ) >> 18)) + B17;
    B19 <= (((32'he9b6c7aa + ((D18&B18) | ((~D18)&C18)) + A18 + w18[ 0 +: 32]) << 20)  |
            ((32'he9b6c7aa + ((D18&B18) | ((~D18)&C18)) + A18 + w18[ 0 +: 32]) >> 12)) + B18;
    B20 <= (((32'hd62f105d + ((D19&B19) | ((~D19)&C19)) + A19                ) <<  5)  |
            ((32'hd62f105d + ((D19&B19) | ((~D19)&C19)) + A19                ) >> 27)) + B19;
    B21 <= (((32'h02441453 + ((D20&B20) | ((~D20)&C20)) + A20                ) <<  9)  |
            ((32'h02441453 + ((D20&B20) | ((~D20)&C20)) + A20                ) >> 23)) + B20;
    B22 <= (((32'hd8a1e681 + ((D21&B21) | ((~D21)&C21)) + A21                ) << 14)  |
            ((32'hd8a1e681 + ((D21&B21) | ((~D21)&C21)) + A21                ) >> 18)) + B21;
    B23 <= (((32'he7d3fbc8 + ((D22&B22) | ((~D22)&C22)) + A22                ) << 20)  |
            ((32'he7d3fbc8 + ((D22&B22) | ((~D22)&C22)) + A22                ) >> 12)) + B22;
    B24 <= (((32'h21e1cde6 + ((D23&B23) | ((~D23)&C23)) + A23                ) <<  5)  |
            ((32'h21e1cde6 + ((D23&B23) | ((~D23)&C23)) + A23                ) >> 27)) + B23;
    B25 <= (((32'hc3370816 + ((D24&B24) | ((~D24)&C24)) + A24                ) <<  9)  |
            ((32'hc3370816 + ((D24&B24) | ((~D24)&C24)) + A24                ) >> 23)) + B24;
    B26 <= (((32'hf4d50d87 + ((D25&B25) | ((~D25)&C25)) + A25                ) << 14)  |
            ((32'hf4d50d87 + ((D25&B25) | ((~D25)&C25)) + A25                ) >> 18)) + B25;
    B27 <= (((32'h455a14ed + ((D26&B26) | ((~D26)&C26)) + A26                ) << 20)  |
            ((32'h455a14ed + ((D26&B26) | ((~D26)&C26)) + A26                ) >> 12)) + B26;
    B28 <= (((32'ha9e3e905 + ((D27&B27) | ((~D27)&C27)) + A27                ) <<  5)  |
            ((32'ha9e3e905 + ((D27&B27) | ((~D27)&C27)) + A27                ) >> 27)) + B27;
    B29 <= (((32'hfcefa478 + ((D28&B28) | ((~D28)&C28)) + A28                ) <<  9)  |
            ((32'hfcefa478 + ((D28&B28) | ((~D28)&C28)) + A28                ) >> 23)) + B28;
    B30 <= (((32'h676f02d9 + ((D29&B29) | ((~D29)&C29)) + A29                ) << 14)  |
            ((32'h676f02d9 + ((D29&B29) | ((~D29)&C29)) + A29                ) >> 18)) + B29;
    B31 <= (((32'h8d2a4c8a + ((D30&B30) | ((~D30)&C30)) + A30                ) << 20)  |
            ((32'h8d2a4c8a + ((D30&B30) | ((~D30)&C30)) + A30                ) >> 12)) + B30;

    B32 <= (((32'hfffa3942 + ( B31  ^   C31   ^   D31 ) + A31                ) <<  4)  |
            ((32'hfffa3942 + ( B31  ^   C31   ^   D31 ) + A31                ) >> 28)) + B31;
    B33 <= (((32'h8771f681 + ( B32  ^   C32   ^   D32 ) + A32                ) << 11)  |
            ((32'h8771f681 + ( B32  ^   C32   ^   D32 ) + A32                ) >> 21)) + B32;
    B34 <= (((32'h6d9d6122 + ( B33  ^   C33   ^   D33 ) + A33                ) << 16)  |
            ((32'h6d9d6122 + ( B33  ^   C33   ^   D33 ) + A33                ) >> 16)) + B33;
    B35 <= (((32'hfde5384c + ( B34  ^   C34   ^   D34 ) + A34                ) << 23)  |
            ((32'hfde5384c + ( B34  ^   C34   ^   D34 ) + A34                ) >>  9)) + B34;
    B36 <= (((32'ha4beea44 + ( B35  ^   C35   ^   D35 ) + A35 + w35[32 +: 32]) <<  4)  |
            ((32'ha4beea44 + ( B35  ^   C35   ^   D35 ) + A35 + w35[32 +: 32]) >> 28)) + B35;
    B37 <= (((32'h4bdecfa9 + ( B36  ^   C36   ^   D36 ) + A36                ) << 11)  |
            ((32'h4bdecfa9 + ( B36  ^   C36   ^   D36 ) + A36                ) >> 21)) + B36;
    B38 <= (((32'hf6bb4b60 + ( B37  ^   C37   ^   D37 ) + A37                ) << 16)  |
            ((32'hf6bb4b60 + ( B37  ^   C37   ^   D37 ) + A37                ) >> 16)) + B37;
    B39 <= (((32'hbebfbc70 + ( B38  ^   C38   ^   D38 ) + A38                ) << 23)  |
            ((32'hbebfbc70 + ( B38  ^   C38   ^   D38 ) + A38                ) >>  9)) + B38;
    B40 <= (((32'h289b7ec6 + ( B39  ^   C39   ^   D39 ) + A39                ) <<  4)  |
            ((32'h289b7ec6 + ( B39  ^   C39   ^   D39 ) + A39                ) >> 28)) + B39;
    B41 <= (((32'heaa127fa + ( B40  ^   C40   ^   D40 ) + A40 + w40[ 0 +: 32]) << 11)  |
            ((32'heaa127fa + ( B40  ^   C40   ^   D40 ) + A40 + w40[ 0 +: 32]) >> 21)) + B40;
    B42 <= (((32'hd4ef3085 + ( B41  ^   C41   ^   D41 ) + A41                ) << 16)  |
            ((32'hd4ef3085 + ( B41  ^   C41   ^   D41 ) + A41                ) >> 16)) + B41;
    B43 <= (((32'h04881d05 + ( B42  ^   C42   ^   D42 ) + A42                ) << 23)  |
            ((32'h04881d05 + ( B42  ^   C42   ^   D42 ) + A42                ) >>  9)) + B42;
    B44 <= (((32'hd9d4d039 + ( B43  ^   C43   ^   D43 ) + A43                ) <<  4)  |
            ((32'hd9d4d039 + ( B43  ^   C43   ^   D43 ) + A43                ) >> 28)) + B43;
    B45 <= (((32'he6db99e5 + ( B44  ^   C44   ^   D44 ) + A44                ) << 11)  |
            ((32'he6db99e5 + ( B44  ^   C44   ^   D44 ) + A44                ) >> 21)) + B44;
    B46 <= (((32'h1fa27cf8 + ( B45  ^   C45   ^   D45 ) + A45                ) << 16)  |
            ((32'h1fa27cf8 + ( B45  ^   C45   ^   D45 ) + A45                ) >> 16)) + B45;
    B47 <= (((32'hc4ac56e5 + ( B46  ^   C46   ^   D46 ) + A46                ) << 23)  |
            ((32'hc4ac56e5 + ( B46  ^   C46   ^   D46 ) + A46                ) >>  9)) + B46;

    B48 <= (((32'hf4292244 + ( C47  ^  (B47   |  ~D47)) + A47 + w47[ 0 +: 32]) <<  6)  |
            ((32'hf4292244 + ( C47  ^  (B47   |  ~D47)) + A47 + w47[ 0 +: 32]) >> 26)) + B47;
    B49 <= (((32'h432aff97 + ( C48  ^  (B48   |  ~D48)) + A48                ) << 10)  |
            ((32'h432aff97 + ( C48  ^  (B48   |  ~D48)) + A48                ) >> 22)) + B48;
    B50 <= (((32'hab9423e7 + ( C49  ^  (B49   |  ~D49)) + A49                ) << 15)  |
            ((32'hab9423e7 + ( C49  ^  (B49   |  ~D49)) + A49                ) >> 17)) + B49;
    B51 <= (((32'hfc93a039 + ( C50  ^  (B50   |  ~D50)) + A50                ) << 21)  |
            ((32'hfc93a039 + ( C50  ^  (B50   |  ~D50)) + A50                ) >> 11)) + B50;
    B52 <= (((32'h655b59c3 + ( C51  ^  (B51   |  ~D51)) + A51                ) <<  6)  |
            ((32'h655b59c3 + ( C51  ^  (B51   |  ~D51)) + A51                ) >> 26)) + B51;
    B53 <= (((32'h8f0ccc92 + ( C52  ^  (B52   |  ~D52)) + A52                ) << 10)  |
            ((32'h8f0ccc92 + ( C52  ^  (B52   |  ~D52)) + A52                ) >> 22)) + B52;
    B54 <= (((32'hffeff47d + ( C53  ^  (B53   |  ~D53)) + A53                ) << 15)  |
            ((32'hffeff47d + ( C53  ^  (B53   |  ~D53)) + A53                ) >> 17)) + B53;
    B55 <= (((32'h85845dd1 + ( C54  ^  (B54   |  ~D54)) + A54 + w54[32 +: 32]) << 21)  |
            ((32'h85845dd1 + ( C54  ^  (B54   |  ~D54)) + A54 + w54[32 +: 32]) >> 11)) + B54;
    B56 <= (((32'h6fa87e4f + ( C55  ^  (B55   |  ~D55)) + A55                ) <<  6)  |
            ((32'h6fa87e4f + ( C55  ^  (B55   |  ~D55)) + A55                ) >> 26)) + B55;
    B57 <= (((32'hfe2ce6e0 + ( C56  ^  (B56   |  ~D56)) + A56                ) << 10)  |
            ((32'hfe2ce6e0 + ( C56  ^  (B56   |  ~D56)) + A56                ) >> 22)) + B56;
    B58 <= (((32'ha3014314 + ( C57  ^  (B57   |  ~D57)) + A57                ) << 15)  |
            ((32'ha3014314 + ( C57  ^  (B57   |  ~D57)) + A57                ) >> 17)) + B57;
    B59 <= (((32'h4e0811a1 + ( C58  ^  (B58   |  ~D58)) + A58                ) << 21)  |
            ((32'h4e0811a1 + ( C58  ^  (B58   |  ~D58)) + A58                ) >> 11)) + B58;
    B60 <= (((32'hf7537e82 + ( C59  ^  (B59   |  ~D59)) + A59                ) <<  6)  |
            ((32'hf7537e82 + ( C59  ^  (B59   |  ~D59)) + A59                ) >> 26)) + B59;
    B61 <= (((32'hbd3af235 + ( C60  ^  (B60   |  ~D60)) + A60                ) << 10)  |
            ((32'hbd3af235 + ( C60  ^  (B60   |  ~D60)) + A60                ) >> 22)) + B60;
    B62 <= (((32'h2ad7d33b + ( C61  ^  (B61   |  ~D61)) + A61                ) << 15)  |
            ((32'h2ad7d33b + ( C61  ^  (B61   |  ~D61)) + A61                ) >> 17)) + B61;
    B63 <= (((32'heb86d391 + ( C62  ^  (B62   |  ~D62)) + A62                ) << 21)  |
            ((32'heb86d391 + ( C62  ^  (B62   |  ~D62)) + A62                ) >> 11)) + B62 + h1;
end

endmodule  // md5